`include "cmos_cells.v"
`include "contador.v"
`include "mux.v"
`include "fifo.v"
`include "referee_1.v"
`include "referee_2.v"
`include "state_machine.v"
`include "demultiplex.v"
`include "multiplexIn.v"
`include "multiplexOut.v"

module tcl();
   // Maquina de Estados
   state_machine maquinaEstados(/*AUTOINST*/
				// Outputs
				.umbral_superior(umbral_superior[2:0]),
				.umbral_inferior(umbral_inferior[2:0]),
				.State		(State[3:0]),
				// Inputs
				.clk		(clk),
				.Umbral_bajo	(Umbral_bajo[2:0]),
				.Umbral_alto	(Umbral_alto[2:0]),
				.reset		(reset),
				.init		(init),
				.empty0		(empty0),
				.empty1		(empty1),
				.empty2		(empty2),
				.empty3		(empty3),
				.empty4		(empty4),
				.empty5		(empty5),
				.empty6		(empty6),
				.empty7		(empty7));
   // Banco Contadores
   mux bancoContadores(/*AUTOINST*/
		       // Outputs
		       .data		(data[4:0]),
		       .valid		(valid),
		       // Inputs
		       .in0		(in0[4:0]),
		       .in1		(in1[4:0]),
		       .in2		(in2[4:0]),
		       .in3		(in3[4:0]),
		       .in4		(in4[4:0]),
		       .state		(state[3:0]),
		       .idx		(idx[2:0]),
		       .req		(req),
		       .clk		(clk));
   // Arbitros
   referee_1 arbitro1(/*AUTOINST*/
		      // Outputs
		      .push_0		(push_0),
		      .push_1		(push_1),
		      .push_2		(push_2),
		      .push_3		(push_3),
		      .pop_0		(pop_0),
		      .pop_1		(pop_1),
		      .pop_2		(pop_2),
		      .pop_3		(pop_3),
		      // Inputs
		      .almost_full_0	(almost_full_0),
		      .almost_full_1	(almost_full_1),
		      .almost_full_2	(almost_full_2),
		      .almost_full_3	(almost_full_3),
		      .empty_0		(empty_0),
		      .empty_1		(empty_1),
		      .empty_2		(empty_2),
		      .empty_3		(empty_3),
		      .clk		(clk),
		      .reset		(reset));
   referee_2 arbitro2(/*AUTOINST*/
		      // Outputs
		      .push_0		(push_0),
		      .push_1		(push_1),
		      .push_2		(push_2),
		      .push_3		(push_3),
		      .pop		(pop),
		      // Inputs
		      .almost_full_0	(almost_full_0),
		      .almost_full_1	(almost_full_1),
		      .almost_full_2	(almost_full_2),
		      .almost_full_3	(almost_full_3),
		      .empty		(empty),
		      .clk		(clk),
		      .reset		(reset));
   // Multiplexor entradas
   multiplexIn multiplexorEntrada(/*AUTOINST*/
				  // Outputs
				  .p0			(p0[11:0]),
				  .p1			(p1[11:0]),
				  .p2			(p2[11:0]),
				  .p3			(p3[11:0]),
				  // Inputs
				  .dataInput		(dataInput[11:0]),
				  .states		(states[3:0]),
				  .clk			(clk));
   // Multiplexor salidas
   multiplexOut multiplexorSalida(/*AUTOINST*/
				  // Outputs
				  .out0			(out0[11:0]),
				  .out1			(out1[11:0]),
				  .out2			(out2[11:0]),
				  .out3			(out3[11:0]),
				  // Inputs
				  .dataInput		(dataInput[11:0]),
				  .states		(states[3:0]),
				  .clk			(clk));
   // Demultiplexor
   demultiplex demultiplexor(/*AUTOINST*/
			     // Outputs
			     .demuxOut		(demuxOut[11:0]),
			     // Inputs
			     .p0		(p0[11:0]),
			     .p1		(p1[11:0]),
			     .p2		(p2[11:0]),
			     .p3		(p3[11:0]),
			     .state		(state[3:0]),
			     .valid0		(valid0),
			     .valid1		(valid1),
			     .valid2		(valid2),
			     .valid3		(valid3),
			     .clk		(clk));
   
   // FIFO Entrada
   fifo fifoIn(/*AUTOINST*/
	       // Outputs
	       .data_out		(data_out[11:0]),
	       .almost_full		(almost_full),
	       .almost_empty		(almost_empty),
	       // Inputs
	       .data_in			(data_in[11:0]),
	       .reset			(reset),
	       .clk			(clk),
	       .umbral_AF_in		(umbral_AF_in[2:0]),
	       .umbral_AE_in		(umbral_AE_in[2:0]),
	       .push			(push),
	       .pop			(pop),
	       .state			(state[3:0]));
   // FIFO Salida
   fifo fifoOut(/*AUTOINST*/
		// Outputs
		.data_out		(data_out[11:0]),
		.almost_full		(almost_full),
		.almost_empty		(almost_empty),
		// Inputs
		.data_in		(data_in[11:0]),
		.reset			(reset),
		.clk			(clk),
		.umbral_AF_in		(umbral_AF_in[2:0]),
		.umbral_AE_in		(umbral_AE_in[2:0]),
		.push			(push),
		.pop			(pop),
		.state			(state[3:0]));
   // Bloque FIFOs entrada
   fifo fifoInP0(/*AUTOINST*/
		 // Outputs
		 .data_out		(data_out[11:0]),
		 .almost_full		(almost_full),
		 .almost_empty		(almost_empty),
		 // Inputs
		 .data_in		(data_in[11:0]),
		 .reset			(reset),
		 .clk			(clk),
		 .umbral_AF_in		(umbral_AF_in[2:0]),
		 .umbral_AE_in		(umbral_AE_in[2:0]),
		 .push			(push),
		 .pop			(pop),
		 .state			(state[3:0]));
   fifo fifoInP1(/*AUTOINST*/
		 // Outputs
		 .data_out		(data_out[11:0]),
		 .almost_full		(almost_full),
		 .almost_empty		(almost_empty),
		 // Inputs
		 .data_in		(data_in[11:0]),
		 .reset			(reset),
		 .clk			(clk),
		 .umbral_AF_in		(umbral_AF_in[2:0]),
		 .umbral_AE_in		(umbral_AE_in[2:0]),
		 .push			(push),
		 .pop			(pop),
		 .state			(state[3:0]));
   fifo fifoInP2(/*AUTOINST*/
		 // Outputs
		 .data_out		(data_out[11:0]),
		 .almost_full		(almost_full),
		 .almost_empty		(almost_empty),
		 // Inputs
		 .data_in		(data_in[11:0]),
		 .reset			(reset),
		 .clk			(clk),
		 .umbral_AF_in		(umbral_AF_in[2:0]),
		 .umbral_AE_in		(umbral_AE_in[2:0]),
		 .push			(push),
		 .pop			(pop),
		 .state			(state[3:0]));
   fifo fifoInP3(/*AUTOINST*/
		 // Outputs
		 .data_out		(data_out[11:0]),
		 .almost_full		(almost_full),
		 .almost_empty		(almost_empty),
		 // Inputs
		 .data_in		(data_in[11:0]),
		 .reset			(reset),
		 .clk			(clk),
		 .umbral_AF_in		(umbral_AF_in[2:0]),
		 .umbral_AE_in		(umbral_AE_in[2:0]),
		 .push			(push),
		 .pop			(pop),
		 .state			(state[3:0]));
   // Bloque FIFOs salida
   fifo fifoOutP0(/*AUTOINST*/
		  // Outputs
		  .data_out		(data_out[11:0]),
		  .almost_full		(almost_full),
		  .almost_empty		(almost_empty),
		  // Inputs
		  .data_in		(data_in[11:0]),
		  .reset		(reset),
		  .clk			(clk),
		  .umbral_AF_in		(umbral_AF_in[2:0]),
		  .umbral_AE_in		(umbral_AE_in[2:0]),
		  .push			(push),
		  .pop			(pop),
		  .state		(state[3:0]));
   fifo fifoOutP1(/*AUTOINST*/
		  // Outputs
		  .data_out		(data_out[11:0]),
		  .almost_full		(almost_full),
		  .almost_empty		(almost_empty),
		  // Inputs
		  .data_in		(data_in[11:0]),
		  .reset		(reset),
		  .clk			(clk),
		  .umbral_AF_in		(umbral_AF_in[2:0]),
		  .umbral_AE_in		(umbral_AE_in[2:0]),
		  .push			(push),
		  .pop			(pop),
		  .state		(state[3:0]));
   fifo fifoOutP2(/*AUTOINST*/
		  // Outputs
		  .data_out		(data_out[11:0]),
		  .almost_full		(almost_full),
		  .almost_empty		(almost_empty),
		  // Inputs
		  .data_in		(data_in[11:0]),
		  .reset		(reset),
		  .clk			(clk),
		  .umbral_AF_in		(umbral_AF_in[2:0]),
		  .umbral_AE_in		(umbral_AE_in[2:0]),
		  .push			(push),
		  .pop			(pop),
		  .state		(state[3:0]));
   fifo fifoOutP3(/*AUTOINST*/
		  // Outputs
		  .data_out		(data_out[11:0]),
		  .almost_full		(almost_full),
		  .almost_empty		(almost_empty),
		  // Inputs
		  .data_in		(data_in[11:0]),
		  .reset		(reset),
		  .clk			(clk),
		  .umbral_AF_in		(umbral_AF_in[2:0]),
		  .umbral_AE_in		(umbral_AE_in[2:0]),
		  .push			(push),
		  .pop			(pop),
		  .state		(state[3:0]));
   
   
endmodule // tcl
