`timescale 	1ns	/ 100ps

`include "cmos_cells.v"
`include "fifo.v"
`include "fifo_str.v"
`include "tester.v"



module testbench;
    
endmodule