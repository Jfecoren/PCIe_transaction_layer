

module tester(
    input [11:0] data_out, data_w,
    input [2:0] addr_w, addr_r,
    input almost_full, almost_empty,
    output reg [11:0] data_in, data_r,
    output reg reset, clk,
    output reg push, pop
);
    
endmodule