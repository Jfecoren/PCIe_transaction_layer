


module fifo(
    
);

endmodule