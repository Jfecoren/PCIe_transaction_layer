

module tester(
    ports
);
    
endmodule